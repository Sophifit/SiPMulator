
library ieee;
use ieee.std_logic_1164.all;

package data_package is

  type s_vector is array(0 to 31) of std_logic_vector(7 downto 0);

end data_package;

package body data_package is

end data_package;